module tb_CSRAM_asyn (
  input clk,    // Clock
  input clk_en, // Clock Enable
  input rst_n,  // Asynchronous reset active low
  
);
CSRAM_asyn CSRAM_asyn_DUT

endmodule